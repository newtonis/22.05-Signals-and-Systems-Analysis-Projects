
module constant_8bit(out);
	output [7:0]out;
	assign out = 24;
	
endmodule