module bit8fixed(out);
	output [7:0]out;
	assign out = 255;
endmodule