module compare_number(a,b);
	input [7:0]a;
	output b;
	assign b = a <= 44;
	
endmodule